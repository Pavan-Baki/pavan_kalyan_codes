vcov merge final.ucdb \
mac_reg_read_test.ucdb \
mac_reg_write_read_test.ucdb \
mac_random_reg_write_read_test.ucdb \
mac_random_reg_wr_nr_test.ucdb \
mac_reg_write_read_reg_model_test.ucdb \
mac_bd_reg_wr_rd_rm_test.ucdb \
mac_reg_rd_rm_test.ucdb \
mac_fd_test.ucdb \
mac_fd_rx_test.ucdb \
mac_fd_tx_rx_test.ucdb \
mac_mii_wctrl_data_tx_test.ucdb \
mac_hd_tx_coll_det_test.ucdb \
mac_fd_tx_pause_frame_test.ucdb

